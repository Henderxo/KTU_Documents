------------------------------------- 

--KTU 2015

--Informatikos fakultetas
--Kompiuteriu katedra
--Kompiuteriu Architektura [P175B125] 
--Kazimieras Bagdonas 

--v1.0

------------------------------------- 
--KTU 2016 

--ditto

--v1.01
--panaikinta "save" mikrokomanda registrams, sutrumpinta ROM eilute nuo 75 iki 69 bitu, nesuderinama su V1.0   

------------------------------------- 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is 
	port (
		RST_ROM 	: in std_logic;
		clk 		: in std_logic;
		ROM_CMD 	: in std_logic_vector(7 downto 0);  
		ROM_Dout 	: out std_logic_vector(1 to 69)
		);
end ROM ;

architecture rtl of ROM is
	
	type memory is array (0 to 255) of std_logic_vector(1 to 69) ; 
	
	constant ROM_CMDln : memory := (  
--                    1         2         3         4         5         6            Dvi komentaro eilutes duoda bitu numerius   
--           123456789012345678901234567890123456789012345678901234567890123456789    (nuo 1 iki 69)
0=>"010000000000000100000000000000000000000000000000000000000000000000000",--Komentarovieta
1=>"010000000000000010000010000000000000000000000000000000000000000000000",--Komentarovieta
2=>"010000000000000001000001000001000000100000000000000000000000000000000",--Komentarovieta
3=>"000000000000000000000000100000000000000000000000000000000000000000000",--Komentarovieta
4=>"000100000000000000000000000000000000000000000000000000000000000000000",--Komentarovieta
5=>"000000001000000000000000000000000000000000000000000100000000000000000",--Komentarovieta
6=>"000010001000000000000000000000000000000000000000000000010000000000000",--Komentarovieta
7=>"0000000010000L0000000000000000000000000000000000001000000000000000000",--Komentarovieta
8=>"001000000000000000000000000000000000000000000000000000000000000000000",--Komentarovieta
9=>"000000000000000000000000000000000000000000010000000000000000000000000",--Komentarovieta
10=>"000001000000000000000000000000000000000000000000000000000010000000000",--Komentarovieta
11=>"000000000000000000000000000000000000000000000000000000000000000000000",--Komentarovieta
12=>"110100000111000000000000000000000000000000000000000000000000000000000",--Komentarovieta
13=>"000000001000000000000000000000000000000000000000001000000000000000000",--Komentarovieta
14=>"000000000000000000000000000000000000000000000000000000000000000000001",--Komentarovieta
15=>"000000000000000000000000000000100000001000000000000000000000000000000",--Komentarovieta
16=>"111010000110000000000000000000000000000000000000000000000000000000000",--Komentarovieta
17=>"001000000000000000000000000000000000000000000000000000000000000000000",--Komentarovieta
18=>"000000000000000000000000000000000000100000000000000000000000000000000",--Komentarovieta
19=>"000000000000000000000000000000000000000000000000000000000010000000000",--Komentarovieta
20=>"000000001000000000000000000000000000000000000000000100000000000000000",--Komentarovieta
21=>"001000000000000000000000000000000000000000000000000000000000000000000",--Komentarovieta
22=>"000000000000000100000000000000000000000000000000000000000000000000000",--Komentarovieta
23=>"000000100000000000000000000000000000000000000000000000000000000000000",--Komentarovieta
24=>"000000001000000000000000000000000000000000000000000100000000000000000",--Komentarovieta
25=>"000000001000000000000000000000000000000000000000000000010000000000000",--Komentarovieta
26=>"001000000000000000000000000000000000000000000000000000000000000000000",--Komentarovieta
27=>"000000000000000000000010000000000000000000000000000010000000000000000",--Komentarovieta
28=>"000000000000000010000001000000000000010000000000000000010000000000000",--Komentarovieta
29=>"000000000000000010000001000000000000010000000000000000000000000000000",--Komentarovieta
30=>"000000000000000010000001000000000000010000000000000000000000000000000",--Komentarovieta
31=>"000000000000000010000001000000000000010000000000000000000000000000000",--Komentarovieta
32=>"000000000000000010000001000000000000010000000000000000000000000000000",--Komentarovieta
33=>"000000000000000010000001000000000000010000000000000000000000000000000",--Komentarovieta
34=>"000000000000000010000001000000000000010000000000000000000000000000000",--Komentarovieta
35=>"000000000000000010000000000000000000000000000000000000000010000000000",--Komentarovieta
36=>"000000000000000000000000000000000000000000000000000000000000000010000",--Komentarovieta
37=>"000000010000000000000000000000000000000000000000000000000000000000000",--Komentarovieta
38=>"000000001000000000000000000000000000000000000000001000000000000000000",--Komentarovieta
39=>"110110010101100000000000000000000000000000000000000000000000000000000",--Komentarovieta
40=>"000000011000000000000000000001000000000000000000000100000000000000000",--Komentarovieta
41=>"000000001000000000000000000000000000000000000000000000010000000000000",--Komentarovieta
42=>"001000000000000000000000000000000000000000010000000000000000000000000",--Komentarovieta
43=>"000010000000000000000000000000000000000000000000000000000000000000000",--Komentarovieta
44=>"000010001000000000000000000000000000000000000000001000000000000000000",--Komentarovieta
45=>"000000000000000000000000000000000000000000000000000000000000000000000",--Komentarovieta
46=>"100010011001100000000000000000000000000000000000000000000000000000000",--Komentarovieta
47=>"000000100000000010000000000000000000000000000000000000000000000000000",--Komentarovieta
48=>"000000101000000000000000000000000000000000000000001000000000000000000",--Komentarovieta
49=>"000000000000000000000000000000000000000000000000000000000000000000000",--Komentarovieta
50=>"111110011010000000000000000000000000000000000000000000000000000000000",--Komentarovieta
51=>"000000000000000000001000000000000000000000000000001000000000000000000",--Komentarovieta
52=>"000000000100000000000000000000000000000000000000000000000000000000000",--Komentarovieta
53=>"000000000000000000000000000000000000000000000000000000000000000000001",--Komentarovieta
54=>"000000000000000000000000000000000000000000000000000000000000000000000",--Komentarovieta
55=>"111010010101100000000000000000000000000000000000000000000000000000000",--Komentarovieta
56=>"101110100010000000000000000000000000000000000000000000000000000000000",--Komentarovieta
57=>"000100000000000000000000000000000000000000000000000000000000000000000",--Komentarovieta
58=>"000000001000000000000000000000000000000000000000000100000000000000000",--Komentarovieta
59=>"000000001000000000000000000000000000000000000000000000010000000000000",--Komentarovieta
60=>"001000000000000100000000000000000000000000000000000000000000000000000",--Komentarovieta
61=>"000100001000000000000000000000000000000000000000000100000000000000000",--Komentarovieta
62=>"000000001000000000000000000000000000000000000000000000010000000000000",--Komentarovieta
63=>"001000000000000100000000000000000000000000000000000000000000000000000",--Komentarovieta
64=>"000000000000000010000000000000000000000000000000000000000000000000000",--Komentarovieta
65=>"000100001000000000000000000000000000000000000000000001000000000000000",--Komentarovieta
66=>"001000000000000100000000000000000000000000000000000000000000000000000",--Komentarovieta
67=>"000000000000000000000100000000000000000000000000000000000000000000000",--Komentarovieta
68=>"000100000000000000000000000000000000000000000000000000000000000000000",--Komentarovieta
69=>"000000000000000000000000000000000000000000000000000000000000000000010",--Komentarovieta

	others => (others => '0') );   
	
	
	
begin
	process (RST_ROM, clk) 
		
	begin
		if RST_ROM'event and RST_ROM = '1' then 
			ROM_Dout <= ROM_CMDln(0);
		elsif clk'event and clk = '0' then
			ROM_Dout <= ROM_CMDln(to_integer(unsigned(ROM_CMD))); 
		end if;
		
	end process;
	
end rtl;